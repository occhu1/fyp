//Receiving FPGA base station by Owen Christopher Chu (26921308)
//This verilog file is used to program the FPGA with the purpose of receiving data from the ADC.
//4 bit lengths are implemented in this module; 7, 11, 15 and 31, but currently only the 7 bit length will be tested. Other bit lengths might be tested in a later date.
//The initial PRBS bit length is 7 bits.
//The push button KEY[3] is used to change the PRBS bit length.
//The push button KEY[2] is used to initiate the DAC when only 1 FPGA is available .
//The 2 left-most 7 segment displays are used to display how many batches of data the board has received from the ADC.
//The PRBS-generated sequence is sent from the ADC interface to the GPIO_1 port.
//The FPGA will generate its own pattern for comparison and error checking.
//LEDR[1:0] will light up if nothing is wrong and LEDR[3:2] will light up if there are errors between the generated pattern and the one received from the ADC.
//LEDR[15:14] will light up if nothing is wrong and LEDR[17:16] will light up if there are errors between the direction connecting between the 2 FPGAs.
module receiver(GPIO_1, GPIO_0, CLOCK_50, KEY, HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7, LEDG, LEDR);
	input 					CLOCK_50;
	input		[3:0]			KEY;
	input		[35:0]		GPIO_1;
	
	output	[35:0]		GPIO_0;
	
	output	[6:0]			HEX0;
	output	[6:0]			HEX1;
	output	[6:0]			HEX2;
	output	[6:0] 		HEX3;
	output	[6:0]			HEX4;
	output	[6:0] 		HEX5;
	output	[6:0] 		HEX6;
	output	[6:0] 		HEX7;
	output	[3:0] 		LEDG;
	output	[17:0] 		LEDR;
	
	reg		[6:0]			prbs07;
	reg		[3:0]			sel_1;				//First digit of the bit length selector
	reg		[3:0]			sel_2;				//Second digit of the bit length selector
	reg						error;
	reg						error2;
	reg						error3;
	reg						error4;
	reg						error5;
	reg		[128:0]		checkin;
	reg		[8:0]			alt_clk;
	reg		[126:0]		preset;
	reg		[126:0]		result;
	reg		[7:0]			buffer0;
	reg		[7:0]			buffer1;
	reg		[7:0]			buffer2;
	reg		[7:0]			buffer3;
	reg		[7:0]			buffer4;
	reg		[7:0]			buffer5;
	reg		[7:0]			buffer6;
	reg		[7:0]			buffer7;
	reg		[7:0]			buffer8;
	reg		[7:0]			buffer9;
	reg		[7:0]			buffer10;
	reg		[7:0]			buffer11;
	reg		[7:0]			buffer12;
	reg		[7:0]			buffer13;
	reg		[7:0]			buffer14;
	reg		[6:0]			buffer15;
	reg						rst_flg;
	reg						rst_flg_old;
	reg		[7:0]			flg_cntr;
	
	//Initial values for the PRBS sequences
	initial prbs07			=		1'b1;
	initial result			=		1'b1;
	initial checkin		= 		1'b1;
	initial sel_1			= 	4'b0000;
	initial sel_2			= 	4'b0111;
	
	integer select			=			0;
	integer old_select	=			0;
	integer error_cntr	=			0;
	integer error_chkr	=			0;
	integer shft_cntr		=			0;
	integer read_cntr		=			0;
	integer position		=			0;
	
	always @ (posedge KEY[3])
	begin
	//Event that occurs when KEY3 is pressed. The current length selector state is saved to old_select and a FSM is implemented to find the next bit length.
	//sel_1 and sel_2 are used to output the bit length value to the 7 segment displays.
	//The selector values 00 represent 7 bits, 01 represent 11 bits, 10 represent 15 bits and 11 represent 31 bits.
	old_select 	= select;
		case(old_select)
		2'b00 : begin
				select =   		1;
				sel_1  = 4'b0001;
				sel_2  = 4'b0001;
			 end
		2'b01 : begin
				select =   		2;
				sel_1  = 4'b0001;
				sel_2  = 4'b0101;
			  end
		2'b10 : begin
				select =   		3;
				sel_1  = 4'b0011;
				sel_2  = 4'b0001;
			  end
		2'b11 : begin
				select =   		0;
				sel_1  = 4'b0000;
				sel_2  = 4'b0111;
			  end
		default : begin
				select =   		0;
				sel_1  = 4'b0001;
				sel_2  = 4'b0111;
			  end
			  endcase
	end
	
	always @(posedge CLOCK_50)
	begin
	//Generates a preset pattern using the same algorithm as the generating FPGA. Checks the received data with the PRBS generated within the board to make sure there were no errors during the transmission of the data.
		alt_clk	= alt_clk + 1'b1;											//Incrementer for other always blocks that require slower clock speeds.
		
		if(shft_cntr < 127)													//Generates a pattern on its own once the board is turned on.
		begin
			preset[shft_cntr] = prbs07[6];
			prbs07 	= {prbs07[5:0] , 	prbs07[6]  ^ prbs07[5]};
			shft_cntr = shft_cntr + 1;
		end
		
		if(read_cntr >= 16)
		begin
		//Transferring all the stored data to the result register once all 16 batches of data has been read. The received data will then be checked against the pattern generated by the board for errors.
			result[7:0]			= buffer0[7:0];
			result[15:8]		= buffer1[7:0];
			result[23:16]		= buffer2[7:0];
			result[31:24]		= buffer3[7:0];
			result[39:32]		= buffer4[7:0];
			result[47:40]		= buffer5[7:0];
			result[55:48]		= buffer6[7:0];
			result[63:56]		= buffer7[7:0];
			result[71:64]		= buffer8[7:0];
			result[79:72]		= buffer9[7:0];
			result[87:80]		= buffer10[7:0];
			result[95:88]		= buffer11[7:0];
			result[103:96]		= buffer12[7:0];
			result[111:104]	= buffer13[7:0];
			result[119:112]	= buffer14[7:0];
			result[126:120]	= buffer15[6:0];
			error					= ~(result == preset);
		end
	end
	
	always @(posedge alt_clk[7])
	begin
	//Data received from the data generating FPGA, used for error checking once all 127 bits of data have been received. 129 bits are stored instead of 127 since a header of 1 followed by a 0 will be sent before the data.
		if(GPIO_1[2] || error_chkr > 0)
		begin
			checkin[error_chkr]	= GPIO_1[2];
			error_chkr				= error_chkr + 1;
		end
		
		if(error_chkr > 129 || error_chkr < 1)
		begin
			error_chkr	= 0;
			error2 		= ~(checkin[128:2] == preset);
		end
	end
	
	always @(posedge GPIO_1[19])
	//Data received from ADC
	begin
		flg_cntr = flg_cntr + 1'b1;
		if(read_cntr >= 16 || rst_flg ^ rst_flg_old)			//Resets the counter used for the switch case below when all 16 batches of data has been read or when the flag reset key has been pressed.
		begin
			read_cntr			= 0;
			flg_cntr				= 0;
			rst_flg_old			= rst_flg;
		end
					
		case(read_cntr)												//As multidimensional arrays can't be implemented, a counter and switch case has been used to store the incoming data to different registers.
		0	:	begin
				buffer0[0]	= GPIO_1[1];
				buffer0[1]	= GPIO_1[3];
				buffer0[2]	= GPIO_1[5];
				buffer0[3]	= GPIO_1[7];
				buffer0[4]	= GPIO_1[9];
				buffer0[5]	= GPIO_1[11];
				buffer0[6]	= GPIO_1[13];
				buffer0[7]	= GPIO_1[15];
				end
		1	:	begin
				buffer1[0]	= GPIO_1[1];
				buffer1[1]	= GPIO_1[3];
				buffer1[2]	= GPIO_1[5];
				buffer1[3]	= GPIO_1[7];
				buffer1[4]	= GPIO_1[9];
				buffer1[5]	= GPIO_1[11];
				buffer1[6]	= GPIO_1[13];
				buffer1[7]	= GPIO_1[15];
				end
		2	:	begin
				buffer2[0]	= GPIO_1[1];
				buffer2[1]	= GPIO_1[3];
				buffer2[2]	= GPIO_1[5];
				buffer2[3]	= GPIO_1[7];
				buffer2[4]	= GPIO_1[9];
				buffer2[5]	= GPIO_1[11];
				buffer2[6]	= GPIO_1[13];
				buffer2[7]	= GPIO_1[15];
				end
		3	:	begin
				buffer3[0]	= GPIO_1[1];
				buffer3[1]	= GPIO_1[3];
				buffer3[2]	= GPIO_1[5];
				buffer3[3]	= GPIO_1[7];
				buffer3[4]	= GPIO_1[9];
				buffer3[5]	= GPIO_1[11];
				buffer3[6]	= GPIO_1[13];
				buffer3[7]	= GPIO_1[15];
				end
		4	:	begin
				buffer4[0]	= GPIO_1[1];
				buffer4[1]	= GPIO_1[3];
				buffer4[2]	= GPIO_1[5];
				buffer4[3]	= GPIO_1[7];
				buffer4[4]	= GPIO_1[9];
				buffer4[5]	= GPIO_1[11];
				buffer4[6]	= GPIO_1[13];
				buffer4[7]	= GPIO_1[15];
				end
		5	:	begin
				buffer5[0]	= GPIO_1[1];
				buffer5[1]	= GPIO_1[3];
				buffer5[2]	= GPIO_1[5];
				buffer5[3]	= GPIO_1[7];
				buffer5[4]	= GPIO_1[9];
				buffer5[5]	= GPIO_1[11];
				buffer5[6]	= GPIO_1[13];
				buffer5[7]	= GPIO_1[15];
				end
		6	:	begin
				buffer6[0]	= GPIO_1[1];
				buffer6[1]	= GPIO_1[3];
				buffer6[2]	= GPIO_1[5];
				buffer6[3]	= GPIO_1[7];
				buffer6[4]	= GPIO_1[9];
				buffer6[5]	= GPIO_1[11];
				buffer6[6]	= GPIO_1[13];
				buffer6[7]	= GPIO_1[15];
				end
		7	:	begin
				buffer7[0]	= GPIO_1[1];
				buffer7[1]	= GPIO_1[3];
				buffer7[2]	= GPIO_1[5];
				buffer7[3]	= GPIO_1[7];
				buffer7[4]	= GPIO_1[9];
				buffer7[5]	= GPIO_1[11];
				buffer7[6]	= GPIO_1[13];
				buffer7[7]	= GPIO_1[15];
				end
		8	:	begin
				buffer8[0]	= GPIO_1[1];
				buffer8[1]	= GPIO_1[3];
				buffer8[2]	= GPIO_1[5];
				buffer8[3]	= GPIO_1[7];
				buffer8[4]	= GPIO_1[9];
				buffer8[5]	= GPIO_1[11];
				buffer8[6]	= GPIO_1[13];
				buffer8[7]	= GPIO_1[15];
				end
		9	:	begin
				buffer9[0]	= GPIO_1[1];
				buffer9[1]	= GPIO_1[3];
				buffer9[2]	= GPIO_1[5];
				buffer9[3]	= GPIO_1[7];
				buffer9[4]	= GPIO_1[9];
				buffer9[5]	= GPIO_1[11];
				buffer9[6]	= GPIO_1[13];
				buffer9[7]	= GPIO_1[15];
				end
		10	:	begin
				buffer10[0]	= GPIO_1[1];
				buffer10[1]	= GPIO_1[3];
				buffer10[2]	= GPIO_1[5];
				buffer10[3]	= GPIO_1[7];
				buffer10[4]	= GPIO_1[9];
				buffer10[5]	= GPIO_1[11];
				buffer10[6]	= GPIO_1[13];
				buffer10[7]	= GPIO_1[15];
				end
		11	:	begin
				buffer11[0]	= GPIO_1[1];
				buffer11[1]	= GPIO_1[3];
				buffer11[2]	= GPIO_1[5];
				buffer11[3]	= GPIO_1[7];
				buffer11[4]	= GPIO_1[9];
				buffer11[5]	= GPIO_1[11];
				buffer11[6]	= GPIO_1[13];
				buffer11[7]	= GPIO_1[15];
				end
		12	:	begin
				buffer12[0]	= GPIO_1[1];
				buffer12[1]	= GPIO_1[3];
				buffer12[2]	= GPIO_1[5];
				buffer12[3]	= GPIO_1[7];
				buffer12[4]	= GPIO_1[9];
				buffer12[5]	= GPIO_1[11];
				buffer12[6]	= GPIO_1[13];
				buffer12[7]	= GPIO_1[15];
				end
		13	:	begin
				buffer13[0]	= GPIO_1[1];
				buffer13[1]	= GPIO_1[3];
				buffer13[2]	= GPIO_1[5];
				buffer13[3]	= GPIO_1[7];
				buffer13[4]	= GPIO_1[9];
				buffer13[5]	= GPIO_1[11];
				buffer13[6]	= GPIO_1[13];
				buffer13[7]	= GPIO_1[15];
				end
		14	:	begin
				buffer14[0]	= GPIO_1[1];
				buffer14[1]	= GPIO_1[3];
				buffer14[2]	= GPIO_1[5];
				buffer14[3]	= GPIO_1[7];
				buffer14[4]	= GPIO_1[9];
				buffer14[5]	= GPIO_1[11];
				buffer14[6]	= GPIO_1[13];
				buffer14[7]	= GPIO_1[15];
				end
		15	:	begin
				buffer15[0]	= GPIO_1[1];
				buffer15[1]	= GPIO_1[3];
				buffer15[2]	= GPIO_1[5];
				buffer15[3]	= GPIO_1[7];
				buffer15[4]	= GPIO_1[9];
				buffer15[5]	= GPIO_1[11];
				buffer15[6]	= GPIO_1[13];
				end
		endcase
		
		read_cntr 				= read_cntr + 1;						//Incrementer to indicate how many batches of data has been read.
	end
	
	always @(posedge KEY[2])
	begin
		rst_flg = rst_flg + 1;											//A toggle to reset the incrementer if the previous read sequence failed and didn't read the exact amount of data batches.
	end
		
	//Reads the result and outputs it to the HEX display	
	hexconverter h1(buffer0[3:0]  , HEX0);
	hexconverter h2(buffer0[7:4]  , HEX1);
	hexconverter h3(buffer1[3:0]  , HEX2);
	hexconverter h4(buffer1[7:4]  , HEX3);
	hexconverter h5(buffer2[3:0]  , HEX4);
	hexconverter h6(buffer2[7:4]  , HEX5);
	hexconverter h7(flg_cntr[3:0]  , HEX6);
	hexconverter h8(flg_cntr[7:4]  , HEX7);
	
	assign LEDG[3:0]  = ~KEY[3:0];
	assign LEDR[0] 	= ~error;
	assign LEDR[1]		= ~error;
	assign LEDR[2]		= error;
	assign LEDR[3]		= error;
	assign LEDR[14]	= ~error2;
	assign LEDR[15]	= ~error2;
	assign LEDR[16]	= error2;
	assign LEDR[17]	= error2;
	assign GPIO_0[1]	=	~KEY[1];										//KEY[1] is used to trigger the DAC if a second FPGA is not available for testing.
endmodule

//Submodule to find the 7-bit values to output to the 7 segment displays.
module hexconverter(digit, hexout);
input [4:0] digit;
output [6:0] hexout;
reg [6:0] hexout;

always @(*)
	case (digit)
	5'b00000 : hexout = 7'b1000000;
	5'b00001 : hexout = 7'b1111001;
	5'b00010 : hexout = 7'b0100100;
	5'b00011 : hexout = 7'b0110000;
	5'b00100 : hexout = 7'b0011001;
	5'b00101 : hexout = 7'b0010010;
	5'b00110 : hexout = 7'b0000010;
	5'b00111 : hexout = 7'b1111000;
	5'b01000 : hexout = 7'b0000000;
	5'b01001 : hexout = 7'b0010000;
	5'b01010 : hexout = 7'b0001000;
	5'b01011 : hexout = 7'b0000011;
	5'b01100 : hexout = 7'b1000110;
	5'b01101 : hexout = 7'b0100001;
	5'b01110 : hexout = 7'b0000110;
	5'b01111 : hexout = 7'b0001110;
	5'b10000 : hexout = 7'b1111111;
	default : hexout = 7'b1111111;
	endcase

endmodule
